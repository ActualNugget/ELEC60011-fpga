
module task1 (
	clk_clk,
	led_pio_external_connection_export);	

	input		clk_clk;
	output	[7:0]	led_pio_external_connection_export;
endmodule
